conectix             k�vbox  Wi2k    �      �  �   ���B��ݮ��O�P����'                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                conectix             k�vbox  Wi2k    �      �  �   ���B��ݮ��O�P����'                                                                                                                                                                                                                                                                                                                                                                                                                                            