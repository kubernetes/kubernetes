conectix             k�qemu  Wi2k    �(     �( �   ���vx{�-�M��*���2                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������conectix             k�qemu  Wi2k    �(     �( �   ���vx{�-�M��*���2                                                                                                                                                                                                                                                                                                                                                                                                                                            