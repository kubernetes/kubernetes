conectix             k�ktap           �      �  �   ���R��rA��+��;�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                tdbatmap      
      ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    conectix             k�ktap           �      �  �   ���R��rA��+��;�                                                                                                                                                                                                                                                                                                                                                                                                                                            